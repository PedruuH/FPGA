library ieee;
use ieee.std_logic_1164.all;
entity minhaFSM is
    port(
        clk, rst, choice : in std_logic;
        output : out std_logic_vector(3 downto 0)
    );
end entity minhaFSM;
architecture arq of minhaFSM is
    type state_type is ( s0, s1, s2, s3 );
    signal current, next_state : state_type;
begin
    process ( clk )
    begin
        if ( clk = '1' ) then
            current <= next_state;
        end if;
    end process;
    process ( current )
    begin
    case current is
        when s0 => 
            output <= "0001";
            if ( rst = '1') then
                next_state <= s1;
            else
                next_state <= s0;
            end if;
        when s1=>
            output <= "0010";
            if ( choice = '1') then
                next_state <= s2;
            else
                next_state <= s3;
            end if;
        when s2=>
            output <= "0100";
            next_state <= s0;
        when s3=>
            output <= "1000";
            next_state <= s0;
        when others =>
            output <= "0000";
            next_state <= s0;
        end case;
    end process;
end architecture arq;